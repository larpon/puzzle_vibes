// Copyright(C) 2022 Lars Pontoppidan. All rights reserved.
// Use of this source code is governed by an MIT license
// that can be found in the LICENSE file.
module main

import shy.lib as shy

const colors = Colors{}

struct Colors {
	blue shy.Color = shy.rgb(24, 143, 216)
}
